----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    13:11:01 11/11/2011 
-- Design Name: 
-- Module Name:    alu - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity alu is
	port(
		op_a, op_b, alu_ops : in   STD_LOGIC_VECTOR (3 downto 0);
		status, result : out  STD_LOGIC_VECTOR (3 downto 0)
	);
end alu;

architecture Behavioral of alu is
  
begin
	process ( op_a, op_b, alu_ops )
		variable carry : std_logic := '0';
		variable zero  : std_logic := '0';
		variable tmp   : unsigned(4 downto 0) := "00000";
  	begin
 
		status <= "0000";
		carry := '0';
		zero := '0';
 
		case alu_ops is
		when "0000" | "0001" => -- add | addc
			tmp := resize(unsigned(op_a), 5) + resize(unsigned(op_b), 5);
			carry := tmp(4);
			result <= std_logic_vector(resize(tmp, result'length));

		when "0010" | "0011" => -- sub | subc
			tmp := resize(unsigned(op_a), 5) - resize(unsigned(op_b), 5);
			carry := tmp(4);
			--if carry = '1' then
			--	tmp := tmp - "00001";
			--end if;
			result <= std_logic_vector(resize(tmp, result'length));

		when "0100" => -- and
			result <= op_a and op_b;

		when "0101" => -- or
			result <= op_a or op_b;

		when "0110" => -- xor
			result <= op_a xor op_b;

		when "0111" => -- cmpa
			result <= not(op_a);

		when others => result <= "1111";
		end case;

		status(2) <= carry;
		if tmp = 0 then
			status(3) <= '1';
		end if;
	end process;

end Behavioral;